formal_tb tb_i (.*);