typedef struct {
    logic [31:0] rs1_val;
    logic [31:0] rs2_val;
} regfile_pkt;
